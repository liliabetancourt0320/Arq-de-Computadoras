//Definir modulo y uss i/o
module _and (input A, input B, output C);
//2. Declrar señales/elementos internos
//NA
//3. Comportamiento del modulo 
	//asignaciones,instancias, conexiones
assign C=A&B;


endmodule;
