module ram_async (
    output reg [7:0] data_out,
    input [7:0] data_in,
    input [7:0] addr,
    input wr, // Se�al de escritura (1 para escribir, 0 para leer)
    input en  // Se�al de habilitaci�n del chip
);

    // Memoria: 256 posiciones de 8 bits cada una
    reg [7:0] memory[0:255];
    
    // Proceso always para gestionar lectura y escritura
    always @* begin
        if (en) begin
            if (wr) begin
                // Operaci�n de escritura:
                // Cuando wr=1 y en=1, se escribe data_in en la direcci�n addr
                memory[addr] = data_in;
                // En la escritura, la salida puede ser indefinida o mantener el �ltimo valor.
                // Aqu� la ponemos en alta impedancia para simular un bus de datos.
                data_out = 8'hZZ; 
            end else begin
                // Operaci�n de lectura:
                // Cuando wr=0 y en=1, se lee el dato de la direcci�n addr
                data_out = memory[addr];
            end
        end else begin
            data_out = 8'hZZ;
        end
    end

endmodule

